127
135
146
159
177
139
150
225
165
197
221
121
195
227
240
155
147
139
204
131
242
230
227
192
240
222
127
162
140
148
142
199
