input(-66) <= "00111011"; --59
input(-65) <= "01011110"; --94
input(-64) <= "00100000"; --32
input(-63) <= "00110111"; --55
input(-62) <= "10011000"; --152
input(-61) <= "01001111"; --79
input(-60) <= "11111000"; --248
input(-59) <= "01101000"; --104
input(-58) <= "00101000"; --40
input(-57) <= "11010111"; --215
input(-56) <= "11010010"; --210
input(-55) <= "11101010"; --234
input(-54) <= "11110011"; --243
input(-53) <= "10011011"; --155
input(-52) <= "10001010"; --138
input(-51) <= "01001101"; --77
input(-50) <= "00110000"; --48
input(-49) <= "00001100"; --12
input(-48) <= "10010000"; --144
input(-47) <= "11010011"; --211
input(-46) <= "00011001"; --25
input(-45) <= "11110110"; --246
input(-44) <= "11110010"; --242
input(-43) <= "01011100"; --92
input(-42) <= "01011011"; --91
input(-41) <= "00011111"; --31
input(-40) <= "11011000"; --216
input(-39) <= "10111111"; --191
input(-38) <= "00100110"; --38
input(-37) <= "00000001"; --1
input(-36) <= "11100111"; --231
input(-35) <= "10000100"; --132
input(-34) <= "11011001"; --217
input(-33) <= "11111100"; --252
input(-32) <= "10010011"; --147
input(-31) <= "00011111"; --31
input(-30) <= "00101100"; --44
input(-29) <= "00011100"; --28
input(-28) <= "01001010"; --74
input(-27) <= "00000011"; --3
input(-26) <= "11001000"; --200
input(-25) <= "11101110"; --238
input(-24) <= "10001011"; --139
input(-23) <= "11010100"; --212
input(-22) <= "11011010"; --218
input(-21) <= "11110100"; --244
input(-20) <= "00010000"; --16
input(-19) <= "10100111"; --167
input(-18) <= "00100010"; --34
input(-17) <= "00110100"; --52
input(-16) <= "01000101"; --69
input(-15) <= "11110101"; --245
input(-14) <= "11011011"; --219
input(-13) <= "10011010"; --154
input(-12) <= "00000010"; --2
input(-11) <= "11010000"; --208
input(-10) <= "10011111"; --159
input(-9) <= "01011110"; --94
input(-8) <= "11011011"; --219
input(-7) <= "01000000"; --64
input(-6) <= "00101010"; --42
input(-5) <= "01111001"; --121
input(-4) <= "01010110"; --86
input(-3) <= "00111100"; --60
input(-2) <= "00100110"; --38
input(-1) <= "00010101"; --21
input(0) <= "11000110"; --198
input(1) <= "11100110"; --230
input(2) <= "10001010"; --138
input(3) <= "00000111"; --7
input(4) <= "11000010"; --194
input(5) <= "01011011"; --91
input(6) <= "00000011"; --3
input(7) <= "10011110"; --158
input(8) <= "00010110"; --22
input(9) <= "00111001"; --57
input(10) <= "11101010"; --234
input(11) <= "01000110"; --70
input(12) <= "00101000"; --40
input(13) <= "01000000"; --64
input(14) <= "01010000"; --80
input(15) <= "10110111"; --183
input(16) <= "10001000"; --136
input(17) <= "00110011"; --51
input(18) <= "11000001"; --193
input(19) <= "01010110"; --86
input(20) <= "10100000"; --160
input(21) <= "10110101"; --181
input(22) <= "01011101"; --93
input(23) <= "11100011"; --227
input(24) <= "11101010"; --234
input(25) <= "11101001"; --233
input(26) <= "01010100"; --84
input(27) <= "01100101"; --101
input(28) <= "00000000"; --0
input(29) <= "10100101"; --165
input(30) <= "10111110"; --190
input(31) <= "00011001"; --25
input(32) <= "01110011"; --115
input(33) <= "01010111"; --87
input(34) <= "11101001"; --233
input(35) <= "00100011"; --35
input(36) <= "11110010"; --242
input(37) <= "11100011"; --227
input(38) <= "11000010"; --194
